module cache_top (
    
);



endmodule : cache_top